//=====================================================================
// Project: 4 core MESI cache design
// File Name: test_lib.svh
// Description: Base test class and list of tests
// Designers: Venky & Suru
//=====================================================================
//TODO: add your testcase files in here
`include "base_test.sv"
`include "Write_hit_read.sv"
`include "write_read_dcache.sv"
`include "write_after_write.sv"
`include "replacement.sv"