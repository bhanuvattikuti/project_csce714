//=====================================================================
// Project: 4 core MESI cache design
// File Name: replacement_write.sv
// Description: Test for read-miss to I-cache
// Designers: Venky & Suru
//=====================================================================

class replacement_write extends base_test;

    //component macro
    `uvm_component_utils(replacement_write)

    //Constructor
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction : new

    //UVM build phase
    function void build_phase(uvm_phase phase);
        uvm_config_wrapper::set(this, "tb.vsequencer.run_phase", "default_sequence", replacement_write_seq::type_id::get());
        super.build_phase(phase);
    endfunction : build_phase

    //UVM run phase()
    task run_phase(uvm_phase phase);
        `uvm_info(get_type_name(), "Executing replacement_write test" , UVM_LOW)
    endtask: run_phase

endclass : replacement_write


// Sequence for a read-miss on I-cache
class replacement_write_seq extends base_vseq;
    //object macro
    `uvm_object_utils(replacement_write_seq)

    cpu_transaction_c trans;

    //constructor
    function new (string name="replacement_write_seq");
        super.new(name);
    endfunction : new

    virtual task body();
    // addr of same set: 4000_000 01 00, 0101, 0110, 0111



        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[1], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC; address == 32'h4001_0000; data==32'h0000_ffff;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[1], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC; address == 32'h4002_0000;data==32'h0000_aaaa;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[1], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC; address == 32'h4003_0000;data==32'h0000_aaaa;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[1], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC; address == 32'h4004_0000;data==32'h0000_aaaa;})
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[1], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC; address == 32'h4005_0000;data==32'h0000_bbbb;})

  `uvm_do_on_with(trans, p_sequencer.cpu_seqr[2], {request_type == READ_REQ; access_cache_type == DCACHE_ACC; address == 32'h4005_0000; })
`uvm_do_on_with(trans, p_sequencer.cpu_seqr[3], {request_type == READ_REQ; access_cache_type == DCACHE_ACC; address == 32'h4001_0000; })


    endtask

endclass : replacement_write_seq
